`default_nettype none

// just a stub to keep the Tiny Tapeout tools happy

module tt_um_example (
    input  wire       Sel_42dB,
    input  wire       Sel_26dB,
    input  wire       vbn,
    input  wire       AGND,
    input  wire       VirGND_FB,
    input  wire       Vin,
    input  wire       Vip,
    output wire       vo,
    output wire       VirGND_Out
);

endmodule
